.title KiCad schematic
U2 NC_01 NC_02 Net-_C3-Pad2_ GND Net-_C1-Pad2_ VSS GND NC_03 NC_04 GND VDD Net-_C1-Pad2_ Net-_C1-Pad2_ Net-_R1-Pad2_ NC_05 NC_06 LM13700
U4 NC_07 NC_08 Net-_C3-Pad2_ Net-_C2-Pad1_ Net-_C2-Pad1_ VSS GND NC_09 NC_10 GND VDD Net-_C3-Pad2_ Net-_C1-Pad2_ GND NC_11 NC_12 LM13700
U3 Net-_C4-Pad1_ NC_13 GND Net-_C2-Pad1_ Net-_C4-Pad1_ VSS GND NC_14 NC_15 NC_16 VDD Net-_C2-Pad1_ GND Net-_C4-Pad1_ NC_17 Net-_C2-Pad1_ LM13700
U7 VSS VDD LM13700
U5 VSS VDD LM13700
U6 VSS VDD LM13700
C4 Net-_C4-Pad1_ GND C
C2 Net-_C2-Pad1_ GND C
C3 GND Net-_C3-Pad2_ C
C1 GND Net-_C1-Pad2_ C
U1 Net-_R1-Pad1_ Net-_R1-Pad2_ Net-_R1-Pad2_ VDD Net-_R1-Pad2_ Net-_R1-Pad2_ LM334M
R1 Net-_R1-Pad1_ Net-_R1-Pad2_ RTRIM
.end
